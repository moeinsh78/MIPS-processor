`timescale 1ns/1ns
module Add32B(input [31:0]A,[31:0]B, output [31:0]S);
  assign S = A + B;
endmodule

